`timescale 1ns/1ns
module muls16 (a,b,y);
    input [15:0] a, b;
    output  [31:0] y;
    wire    [15:0] ab0 = a & {16{b[0]}};
    wire    [15:0] ab1 = a & {16{b[1]}};
    wire    [15:0] ab2 = a & {16{b[2]}};
    wire    [15:0] ab3 = a & {16{b[3]}};
    wire    [15:0] ab4 = a & {16{b[4]}};
    wire    [15:0] ab5 = a & {16{b[5]}};
    wire    [15:0] ab6 = a & {16{b[6]}};
    wire    [15:0] ab7 = a & {16{b[7]}};
    wire    [15:0] ab8 = a & {16{b[8]}};
    wire    [15:0] ab9 = a & {16{b[9]}};
    wire    [15:0] ab10 = a & {16{b[10]}};
    wire    [15:0] ab11 = a & {16{b[11]}};
    wire    [15:0] ab12 = a & {16{b[12]}};
    wire    [15:0] ab13 = a & {16{b[13]}};
    wire    [15:0] ab14 = a & {16{b[14]}};
    wire    [15:0] ab15 = a & {16{b[15]}};

    // Serial Adder
    // Yi has 32 terms
    assign y = ({16'b1, ~ab0[15], ab0[14:0]}
               +{15'b0, ~ab1[15], ab1[14:0],1'b0}
               +{14'b0, ~ab2[15], ab2[14:0],2'b0}
               +{13'b0, ~ab3[15], ab3[14:0],3'b0}
               +{12'b0, ~ab4[15], ab4[14:0],4'b0}
               +{11'b0, ~ab5[15], ab5[14:0],5'b0}
               +{10'b0, ~ab6[15], ab6[14:0],6'b0}
               +{9'b0,  ~ab7[15], ab7[14:0],7'b0}
                 +{8'b0,~ab8[15], ab8[14:0],8'b0}
                +{7'b0, ~ab9[15], ab9[14:0],9'b0}
               +{6'b0, ~ab10[15], ab10[14:0],10'b0}
               +{5'b0, ~ab11[15], ab11[14:0],11'b0}
                +{4'b0,~ab12[15], ab12[14:0],12'b0}
              + {3'b0, ~ab13[15], ab13[14:0],13'b0}
               +{2'b0, ~ab14[15], ab14[14:0],14'b0}
               + {1'b1, ab15[15],~ab15[14:0],15'b0});
   // Parallel Adder
   // Yi has i+1 terms (i starting from bottom).
    /* assign y = {1, */
    /*                                                                                                                                    ab15[15], */
    /*                                                                                                                         ~ab14[15]+~ab15[14], */
    /*                                                                                                                ab13[15]+ab14[14]+~ab15[13], */
    /*                                                                                                       ~ab12[15]+ab13[14]+ab14[13]+~ab15[12], */
    /*                                                                                              ~ab11[15]+ab12[14]+ab13[13]+ab14[12]+~ab15[11], */
    /*                                                                                     ~ab10[15]+ab11[14]+ab12[13]+ab13[12]+ab14[11]+~ab15[10], */
    /*                                                                             ~ab9[15]+ab10[14]+ab11[13]+ab12[12]+ab13[11]+ab14[10]+~ab15[9], */
    /*                                                                     ~ab8[15]+ab9[14]+ab10[13]+ab11[12]+ab12[11]+ab13[10]+ab14[9]+~ab15[8], */
    /*                                                             ~ab7[15]+ab8[14]+ab9[13]+ab10[12]+ab11[11]+ab12[10]+ab13[9]+ab14[8]+~ab15[7], */
    /*                                                     ~ab6[15]+ab7[14]+ab8[13]+ab9[12]+ab10[11]+ab11[10]+ab12[9]+ab13[8]+ab14[7]+~ab15[6], */
    /*                                             ~ab5[15]+ab6[14]+ab7[13]+ab8[12]+ab9[11]+ab10[10]+ab11[9]+ab12[8]+ab13[7]+ab14[6]+~ab15[5], */
    /*                                     ~ab4[15]+ab5[14]+ab6[13]+ab7[12]+ab8[11]+ab9[10]+ab10[9]+ab11[8]+ab12[7]+ab13[6]+ab14[5]+~ab15[4], */
    /*                             ~ab3[15]+ab4[14]+ab5[13]+ab6[12]+ab7[11]+ab8[10]+ab9[9]+ab10[8]+ab11[7]+ab12[6]+ab13[5]+ab14[4]+~ab15[3], */
    /*                     ~ab2[15]+ab3[14]+ab4[13]+ab5[12]+ab6[11]+ab7[10]+ab8[9]+ab9[8]+ab10[7]+ab11[6]+ab12[5]+ab13[4]+ab14[3]+~ab15[2], */
    /*           1+~ab1[15]+ab2[14]+ab3[13]+ab4[12]+ab5[11]+ab6[10]+ab7[9]+ab8[8]+ab9[7]+ab10[6]+ab11[5]+ab12[4]+ab13[3]+ab14[2]+~ab15[1], */
    /*     ~ab0[15]+ab1[14]+ab2[13]+ab3[12]+ab4[11]+ab5[10]+ab6[9]+ab7[8]+ab8[7]+ab9[6]+ab10[5]+ab11[4]+ab12[3]+ab13[2]+ab14[1]+~ab15[0], */
    /*     ab0[14]+ab1[13]+ab2[12]+ab3[11]+ab4[10]+ab5[9]+ab6[8]+ab7[7]+ab8[6]+ab9[5]+ab10[4]+ab11[3]+ab12[2]+ab13[1]+ab14[0], */
    /*     ab0[13]+ab1[12]+ab2[11]+ab3[10]+ab4[9]+ab5[8]+ab6[7]+ab7[6]+ab8[5]+ab9[4]+ab10[3]+ab11[2]+ab12[1]+ab13[0], */
    /*     ab0[12]+ab1[11]+ab2[10]+ab3[9]+ab4[8]+ab5[7]+ab6[6]+ab7[5]+ab8[4]+ab9[3]+ab10[2]+ab11[1]+ab12[0], */
    /*     ab0[11]+ab1[10]+ab2[9]+ab3[8]+ab4[7]+ab5[6]+ab6[5]+ab7[4]+ab8[3]+ab9[2]+ab10[1]+ab11[0], */
    /*     ab0[10]+ab1[9]+ab2[8]+ab3[7]+ab4[6]+ab5[5]+ab6[4]+ab7[3]+ab8[2]+ab9[1]+ab10[0], */
    /*     ab0[9]+ab1[8]+ab2[7]+ab3[6]+ab4[5]+ab5[4]+ab6[3]+ab7[2]+ab8[1]+ab9[0], */
    /*     ab0[8]+ab1[7]+ab2[6]+ab3[5]+ab4[4]+ab5[3]+ab6[2]+ab7[1]+ab8[0], */
    /*     ab0[7]+ab1[6]+ab2[5]+ab3[4]+ab4[3]+ab5[2]+ab6[1]+ab7[0], */
    /*     ab0[6]+ab1[5]+ab2[4]+ab3[3]+ab4[2]+ab5[1]+ab6[0], */
    /*     ab0[5]+ab1[4]+ab2[3]+ab3[2]+ab4[1]+ab5[0], */
    /*     ab0[4]+ab1[3]+ab2[2]+ab3[1]+ab4[0], */
    /*     ab0[3]+ab1[2]+ab2[1]+ab3[0], */
    /*     ab0[2]+ab1[1]+ab2[0], */
    /*     ab0[1]+ab1[0], */
    /*     ab0[0] */
    /* }; */
endmodule
